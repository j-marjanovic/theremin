///////////////////////////////////////////////////////////////////////////////
//   __  __          _____      _         _   _  ______      _______ _____   //
//  |  \/  |   /\   |  __ \    | |  /\   | \ | |/ __ \ \    / /_   _/ ____|  //
//  | \  / |  /  \  | |__) |   | | /  \  |  \| | |  | \ \  / /  | || |       //
//  | |\/| | / /\ \ |  _  /_   | |/ /\ \ | . ` | |  | |\ \/ /   | || |       //
//  | |  | |/ ____ \| | \ \ |__| / ____ \| |\  | |__| | \  /   _| || |____   //
//  |_|  |_/_/    \_\_|  \_\____/_/    \_\_| \_|\____/   \/   |_____\_____|  //
//                                                                           //
//                          JAN MARJANOVIC, 2014                             //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////


module delay # (
	parameter SIG_BITS	= 16,
	parameter BLEND_B	= 10,	
	parameter DLY_B		= 14,
	parameter FDB_B		= 10
)(
	//------------ Clk and reset ------------
	input 						clk,
	input						reset_n,
	//------------ Input --------------------
	input		[SIG_BITS-1:0]	in,
	//------------ Output -------------------
	output logic [SIG_BITS-1:0]	out,
	//------------ Control ------------------
	input		[BLEND_B-1:0]	blend,
	input		[DLY_B-1:0]		delay,
	input		[FDB_B-1:0]		feedbk	
);




endmodule
