///////////////////////////////////////////////////////////////////////////////
//   __  __          _____      _         _   _  ______      _______ _____   //
//  |  \/  |   /\   |  __ \    | |  /\   | \ | |/ __ \ \    / /_   _/ ____|  //
//  | \  / |  /  \  | |__) |   | | /  \  |  \| | |  | \ \  / /  | || |       //
//  | |\/| | / /\ \ |  _  /_   | |/ /\ \ | . ` | |  | |\ \/ /   | || |       //
//  | |  | |/ ____ \| | \ \ |__| / ____ \| |\  | |__| | \  /   _| || |____   //
//  |_|  |_/_/    \_\_|  \_\____/_/    \_\_| \_|\____/   \/   |_____\_____|  //
//                                                                           //
//                          JAN MARJANOVIC, 2014                             //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////


module tone_gen # (
	parameter F_BITS	= 12,
	parameter A_BITS	= 3,
	parameter SIG_BITS	= 16
)(
	//------------ Clk and reset ------------
	input 						clk,
	input						reset_n,
	//------------ Input --------------------
	input		[F_BITS-1:0]	freq,
	//------------ Tone Control -------------
	input		[A_BITS-1:0]	a16,
	input		[A_BITS-1:0]	a8,
	input		[A_BITS-1:0]	a5,
	input		[A_BITS-1:0]	a4,
	//------------ Output control -----------
	output reg	[SIG_BITS-1:0]	out
);


endmodule
