

module mem_qsys_top;

mem_controller_tb mem_controller_tb_inst();
mem_qsys_program mem_qsys_program_inst();


endmodule
