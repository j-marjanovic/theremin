///////////////////////////////////////////////////////////////////////////////
//   __  __          _____      _         _   _  ______      _______ _____   //
//  |  \/  |   /\   |  __ \    | |  /\   | \ | |/ __ \ \    / /_   _/ ____|  //
//  | \  / |  /  \  | |__) |   | | /  \  |  \| | |  | \ \  / /  | || |       //
//  | |\/| | / /\ \ |  _  /_   | |/ /\ \ | . ` | |  | |\ \/ /   | || |       //
//  | |  | |/ ____ \| | \ \ |__| / ____ \| |\  | |__| | \  /   _| || |____   //
//  |_|  |_/_/    \_\_|  \_\____/_/    \_\_| \_|\____/   \/   |_____\_____|  //
//                                                                           //
//                          JAN MARJANOVIC, 2014                             //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////
//                                                                           //
//  out = (a * mix + b * (2**M_WIDTH - mix) ) / 2**M_WIDTH                   //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////

module mixer #(
	parameter D_WIDTH 	= 16,
	parameter M_WIDTH 	= 4
)(
	input  [D_WIDTH-1:0] 	a,
	input  [D_WIDTH-1:0] 	b,
	input  [M_WIDTH-1:0] 	mix,
	output [D_WIDTH-1:0]	out
);

wire [M_WIDTH-1:0] antimix = 2**M_WIDTH - 1 - mix;

wire [D_WIDTH+M_WIDTH:0] out_full = (mix*a) + (antimix*b);

assign out = out_full[D_WIDTH+M_WIDTH:M_WIDTH];


endmodule

//=============================================================================
module mixer_tb;

logic [15:0] a, b;
logic [3:0]  mix;
wire  [15:0] out;

mixer mixer_inst( .* );


initial begin
	mix = 0;
	a	= 0;
	b	= 0;
	#1;

	b 	= 100;
	#1;

	b	= 15000;
	#1;

	a	= 15000;
	#1;

	mix	= 5;
	#1;

	mix = 4'b1111;
	#1;

	b	= 0;
	#1;
	
	
	a	= 100;
	#1;

	a	= 1000;
	b	= 100;
	#1;

	for(int i = 0; i < 16; i++) begin
		mix = i;
		#1;
	end
	
	

end


endmodule
