
initial begin
    LUT_sin[0] = 16'd32768;
    LUT_sin[1] = 16'd33170;
    LUT_sin[2] = 16'd33572;
    LUT_sin[3] = 16'd33974;
    LUT_sin[4] = 16'd34375;
    LUT_sin[5] = 16'd34777;
    LUT_sin[6] = 16'd35178;
    LUT_sin[7] = 16'd35579;
    LUT_sin[8] = 16'd35979;
    LUT_sin[9] = 16'd36379;
    LUT_sin[10] = 16'd36779;
    LUT_sin[11] = 16'd37177;
    LUT_sin[12] = 16'd37575;
    LUT_sin[13] = 16'd37973;
    LUT_sin[14] = 16'd38369;
    LUT_sin[15] = 16'd38765;
    LUT_sin[16] = 16'd39160;
    LUT_sin[17] = 16'd39554;
    LUT_sin[18] = 16'd39947;
    LUT_sin[19] = 16'd40339;
    LUT_sin[20] = 16'd40729;
    LUT_sin[21] = 16'd41119;
    LUT_sin[22] = 16'd41507;
    LUT_sin[23] = 16'd41894;
    LUT_sin[24] = 16'd42279;
    LUT_sin[25] = 16'd42663;
    LUT_sin[26] = 16'd43046;
    LUT_sin[27] = 16'd43427;
    LUT_sin[28] = 16'd43806;
    LUT_sin[29] = 16'd44184;
    LUT_sin[30] = 16'd44560;
    LUT_sin[31] = 16'd44934;
    LUT_sin[32] = 16'd45307;
    LUT_sin[33] = 16'd45677;
    LUT_sin[34] = 16'd46046;
    LUT_sin[35] = 16'd46413;
    LUT_sin[36] = 16'd46777;
    LUT_sin[37] = 16'd47140;
    LUT_sin[38] = 16'd47500;
    LUT_sin[39] = 16'd47858;
    LUT_sin[40] = 16'd48214;
    LUT_sin[41] = 16'd48567;
    LUT_sin[42] = 16'd48918;
    LUT_sin[43] = 16'd49267;
    LUT_sin[44] = 16'd49613;
    LUT_sin[45] = 16'd49957;
    LUT_sin[46] = 16'd50298;
    LUT_sin[47] = 16'd50636;
    LUT_sin[48] = 16'd50972;
    LUT_sin[49] = 16'd51305;
    LUT_sin[50] = 16'd51635;
    LUT_sin[51] = 16'd51962;
    LUT_sin[52] = 16'd52287;
    LUT_sin[53] = 16'd52608;
    LUT_sin[54] = 16'd52927;
    LUT_sin[55] = 16'd53242;
    LUT_sin[56] = 16'd53555;
    LUT_sin[57] = 16'd53864;
    LUT_sin[58] = 16'd54170;
    LUT_sin[59] = 16'd54473;
    LUT_sin[60] = 16'd54772;
    LUT_sin[61] = 16'd55069;
    LUT_sin[62] = 16'd55362;
    LUT_sin[63] = 16'd55651;
    LUT_sin[64] = 16'd55937;
    LUT_sin[65] = 16'd56220;
    LUT_sin[66] = 16'd56499;
    LUT_sin[67] = 16'd56774;
    LUT_sin[68] = 16'd57046;
    LUT_sin[69] = 16'd57314;
    LUT_sin[70] = 16'd57579;
    LUT_sin[71] = 16'd57840;
    LUT_sin[72] = 16'd58097;
    LUT_sin[73] = 16'd58350;
    LUT_sin[74] = 16'd58599;
    LUT_sin[75] = 16'd58845;
    LUT_sin[76] = 16'd59086;
    LUT_sin[77] = 16'd59324;
    LUT_sin[78] = 16'd59557;
    LUT_sin[79] = 16'd59787;
    LUT_sin[80] = 16'd60012;
    LUT_sin[81] = 16'd60234;
    LUT_sin[82] = 16'd60451;
    LUT_sin[83] = 16'd60664;
    LUT_sin[84] = 16'd60873;
    LUT_sin[85] = 16'd61077;
    LUT_sin[86] = 16'd61278;
    LUT_sin[87] = 16'd61474;
    LUT_sin[88] = 16'd61665;
    LUT_sin[89] = 16'd61853;
    LUT_sin[90] = 16'd62036;
    LUT_sin[91] = 16'd62214;
    LUT_sin[92] = 16'd62389;
    LUT_sin[93] = 16'd62558;
    LUT_sin[94] = 16'd62723;
    LUT_sin[95] = 16'd62884;
    LUT_sin[96] = 16'd63040;
    LUT_sin[97] = 16'd63192;
    LUT_sin[98] = 16'd63339;
    LUT_sin[99] = 16'd63481;
    LUT_sin[100] = 16'd63619;
    LUT_sin[101] = 16'd63752;
    LUT_sin[102] = 16'd63881;
    LUT_sin[103] = 16'd64004;
    LUT_sin[104] = 16'd64124;
    LUT_sin[105] = 16'd64238;
    LUT_sin[106] = 16'd64348;
    LUT_sin[107] = 16'd64452;
    LUT_sin[108] = 16'd64553;
    LUT_sin[109] = 16'd64648;
    LUT_sin[110] = 16'd64738;
    LUT_sin[111] = 16'd64824;
    LUT_sin[112] = 16'd64905;
    LUT_sin[113] = 16'd64981;
    LUT_sin[114] = 16'd65052;
    LUT_sin[115] = 16'd65118;
    LUT_sin[116] = 16'd65180;
    LUT_sin[117] = 16'd65236;
    LUT_sin[118] = 16'd65288;
    LUT_sin[119] = 16'd65335;
    LUT_sin[120] = 16'd65377;
    LUT_sin[121] = 16'd65414;
    LUT_sin[122] = 16'd65446;
    LUT_sin[123] = 16'd65473;
    LUT_sin[124] = 16'd65495;
    LUT_sin[125] = 16'd65512;
    LUT_sin[126] = 16'd65525;
    LUT_sin[127] = 16'd65532;
    LUT_sin[128] = 16'd65535;
    LUT_sin[129] = 16'd65532;
    LUT_sin[130] = 16'd65525;
    LUT_sin[131] = 16'd65512;
    LUT_sin[132] = 16'd65495;
    LUT_sin[133] = 16'd65473;
    LUT_sin[134] = 16'd65446;
    LUT_sin[135] = 16'd65414;
    LUT_sin[136] = 16'd65377;
    LUT_sin[137] = 16'd65335;
    LUT_sin[138] = 16'd65288;
    LUT_sin[139] = 16'd65236;
    LUT_sin[140] = 16'd65180;
    LUT_sin[141] = 16'd65118;
    LUT_sin[142] = 16'd65052;
    LUT_sin[143] = 16'd64981;
    LUT_sin[144] = 16'd64905;
    LUT_sin[145] = 16'd64824;
    LUT_sin[146] = 16'd64738;
    LUT_sin[147] = 16'd64648;
    LUT_sin[148] = 16'd64553;
    LUT_sin[149] = 16'd64452;
    LUT_sin[150] = 16'd64348;
    LUT_sin[151] = 16'd64238;
    LUT_sin[152] = 16'd64124;
    LUT_sin[153] = 16'd64004;
    LUT_sin[154] = 16'd63881;
    LUT_sin[155] = 16'd63752;
    LUT_sin[156] = 16'd63619;
    LUT_sin[157] = 16'd63481;
    LUT_sin[158] = 16'd63339;
    LUT_sin[159] = 16'd63192;
    LUT_sin[160] = 16'd63040;
    LUT_sin[161] = 16'd62884;
    LUT_sin[162] = 16'd62723;
    LUT_sin[163] = 16'd62558;
    LUT_sin[164] = 16'd62389;
    LUT_sin[165] = 16'd62214;
    LUT_sin[166] = 16'd62036;
    LUT_sin[167] = 16'd61853;
    LUT_sin[168] = 16'd61665;
    LUT_sin[169] = 16'd61474;
    LUT_sin[170] = 16'd61278;
    LUT_sin[171] = 16'd61077;
    LUT_sin[172] = 16'd60873;
    LUT_sin[173] = 16'd60664;
    LUT_sin[174] = 16'd60451;
    LUT_sin[175] = 16'd60234;
    LUT_sin[176] = 16'd60012;
    LUT_sin[177] = 16'd59787;
    LUT_sin[178] = 16'd59557;
    LUT_sin[179] = 16'd59324;
    LUT_sin[180] = 16'd59086;
    LUT_sin[181] = 16'd58845;
    LUT_sin[182] = 16'd58599;
    LUT_sin[183] = 16'd58350;
    LUT_sin[184] = 16'd58097;
    LUT_sin[185] = 16'd57840;
    LUT_sin[186] = 16'd57579;
    LUT_sin[187] = 16'd57314;
    LUT_sin[188] = 16'd57046;
    LUT_sin[189] = 16'd56774;
    LUT_sin[190] = 16'd56499;
    LUT_sin[191] = 16'd56220;
    LUT_sin[192] = 16'd55937;
    LUT_sin[193] = 16'd55651;
    LUT_sin[194] = 16'd55362;
    LUT_sin[195] = 16'd55069;
    LUT_sin[196] = 16'd54772;
    LUT_sin[197] = 16'd54473;
    LUT_sin[198] = 16'd54170;
    LUT_sin[199] = 16'd53864;
    LUT_sin[200] = 16'd53555;
    LUT_sin[201] = 16'd53242;
    LUT_sin[202] = 16'd52927;
    LUT_sin[203] = 16'd52608;
    LUT_sin[204] = 16'd52287;
    LUT_sin[205] = 16'd51962;
    LUT_sin[206] = 16'd51635;
    LUT_sin[207] = 16'd51305;
    LUT_sin[208] = 16'd50972;
    LUT_sin[209] = 16'd50636;
    LUT_sin[210] = 16'd50298;
    LUT_sin[211] = 16'd49957;
    LUT_sin[212] = 16'd49613;
    LUT_sin[213] = 16'd49267;
    LUT_sin[214] = 16'd48918;
    LUT_sin[215] = 16'd48567;
    LUT_sin[216] = 16'd48214;
    LUT_sin[217] = 16'd47858;
    LUT_sin[218] = 16'd47500;
    LUT_sin[219] = 16'd47140;
    LUT_sin[220] = 16'd46777;
    LUT_sin[221] = 16'd46413;
    LUT_sin[222] = 16'd46046;
    LUT_sin[223] = 16'd45677;
    LUT_sin[224] = 16'd45307;
    LUT_sin[225] = 16'd44934;
    LUT_sin[226] = 16'd44560;
    LUT_sin[227] = 16'd44184;
    LUT_sin[228] = 16'd43806;
    LUT_sin[229] = 16'd43427;
    LUT_sin[230] = 16'd43046;
    LUT_sin[231] = 16'd42663;
    LUT_sin[232] = 16'd42279;
    LUT_sin[233] = 16'd41894;
    LUT_sin[234] = 16'd41507;
    LUT_sin[235] = 16'd41119;
    LUT_sin[236] = 16'd40729;
    LUT_sin[237] = 16'd40339;
    LUT_sin[238] = 16'd39947;
    LUT_sin[239] = 16'd39554;
    LUT_sin[240] = 16'd39160;
    LUT_sin[241] = 16'd38765;
    LUT_sin[242] = 16'd38369;
    LUT_sin[243] = 16'd37973;
    LUT_sin[244] = 16'd37575;
    LUT_sin[245] = 16'd37177;
    LUT_sin[246] = 16'd36779;
    LUT_sin[247] = 16'd36379;
    LUT_sin[248] = 16'd35979;
    LUT_sin[249] = 16'd35579;
    LUT_sin[250] = 16'd35178;
    LUT_sin[251] = 16'd34777;
    LUT_sin[252] = 16'd34375;
    LUT_sin[253] = 16'd33974;
    LUT_sin[254] = 16'd33572;
    LUT_sin[255] = 16'd33170;
    LUT_sin[256] = 16'd32768;
    LUT_sin[257] = 16'd32365;
    LUT_sin[258] = 16'd31963;
    LUT_sin[259] = 16'd31561;
    LUT_sin[260] = 16'd31160;
    LUT_sin[261] = 16'd30758;
    LUT_sin[262] = 16'd30357;
    LUT_sin[263] = 16'd29956;
    LUT_sin[264] = 16'd29556;
    LUT_sin[265] = 16'd29156;
    LUT_sin[266] = 16'd28756;
    LUT_sin[267] = 16'd28358;
    LUT_sin[268] = 16'd27960;
    LUT_sin[269] = 16'd27562;
    LUT_sin[270] = 16'd27166;
    LUT_sin[271] = 16'd26770;
    LUT_sin[272] = 16'd26375;
    LUT_sin[273] = 16'd25981;
    LUT_sin[274] = 16'd25588;
    LUT_sin[275] = 16'd25196;
    LUT_sin[276] = 16'd24806;
    LUT_sin[277] = 16'd24416;
    LUT_sin[278] = 16'd24028;
    LUT_sin[279] = 16'd23641;
    LUT_sin[280] = 16'd23256;
    LUT_sin[281] = 16'd22872;
    LUT_sin[282] = 16'd22489;
    LUT_sin[283] = 16'd22108;
    LUT_sin[284] = 16'd21729;
    LUT_sin[285] = 16'd21351;
    LUT_sin[286] = 16'd20975;
    LUT_sin[287] = 16'd20601;
    LUT_sin[288] = 16'd20228;
    LUT_sin[289] = 16'd19858;
    LUT_sin[290] = 16'd19489;
    LUT_sin[291] = 16'd19122;
    LUT_sin[292] = 16'd18758;
    LUT_sin[293] = 16'd18395;
    LUT_sin[294] = 16'd18035;
    LUT_sin[295] = 16'd17677;
    LUT_sin[296] = 16'd17321;
    LUT_sin[297] = 16'd16968;
    LUT_sin[298] = 16'd16617;
    LUT_sin[299] = 16'd16268;
    LUT_sin[300] = 16'd15922;
    LUT_sin[301] = 16'd15578;
    LUT_sin[302] = 16'd15237;
    LUT_sin[303] = 16'd14899;
    LUT_sin[304] = 16'd14563;
    LUT_sin[305] = 16'd14230;
    LUT_sin[306] = 16'd13900;
    LUT_sin[307] = 16'd13573;
    LUT_sin[308] = 16'd13248;
    LUT_sin[309] = 16'd12927;
    LUT_sin[310] = 16'd12608;
    LUT_sin[311] = 16'd12293;
    LUT_sin[312] = 16'd11980;
    LUT_sin[313] = 16'd11671;
    LUT_sin[314] = 16'd11365;
    LUT_sin[315] = 16'd11062;
    LUT_sin[316] = 16'd10763;
    LUT_sin[317] = 16'd10466;
    LUT_sin[318] = 16'd10173;
    LUT_sin[319] = 16'd9884;
    LUT_sin[320] = 16'd9598;
    LUT_sin[321] = 16'd9315;
    LUT_sin[322] = 16'd9036;
    LUT_sin[323] = 16'd8761;
    LUT_sin[324] = 16'd8489;
    LUT_sin[325] = 16'd8221;
    LUT_sin[326] = 16'd7956;
    LUT_sin[327] = 16'd7695;
    LUT_sin[328] = 16'd7438;
    LUT_sin[329] = 16'd7185;
    LUT_sin[330] = 16'd6936;
    LUT_sin[331] = 16'd6690;
    LUT_sin[332] = 16'd6449;
    LUT_sin[333] = 16'd6211;
    LUT_sin[334] = 16'd5978;
    LUT_sin[335] = 16'd5748;
    LUT_sin[336] = 16'd5523;
    LUT_sin[337] = 16'd5301;
    LUT_sin[338] = 16'd5084;
    LUT_sin[339] = 16'd4871;
    LUT_sin[340] = 16'd4662;
    LUT_sin[341] = 16'd4458;
    LUT_sin[342] = 16'd4257;
    LUT_sin[343] = 16'd4061;
    LUT_sin[344] = 16'd3870;
    LUT_sin[345] = 16'd3682;
    LUT_sin[346] = 16'd3499;
    LUT_sin[347] = 16'd3321;
    LUT_sin[348] = 16'd3146;
    LUT_sin[349] = 16'd2977;
    LUT_sin[350] = 16'd2812;
    LUT_sin[351] = 16'd2651;
    LUT_sin[352] = 16'd2495;
    LUT_sin[353] = 16'd2343;
    LUT_sin[354] = 16'd2196;
    LUT_sin[355] = 16'd2054;
    LUT_sin[356] = 16'd1916;
    LUT_sin[357] = 16'd1783;
    LUT_sin[358] = 16'd1654;
    LUT_sin[359] = 16'd1531;
    LUT_sin[360] = 16'd1411;
    LUT_sin[361] = 16'd1297;
    LUT_sin[362] = 16'd1187;
    LUT_sin[363] = 16'd1083;
    LUT_sin[364] = 16'd982;
    LUT_sin[365] = 16'd887;
    LUT_sin[366] = 16'd797;
    LUT_sin[367] = 16'd711;
    LUT_sin[368] = 16'd630;
    LUT_sin[369] = 16'd554;
    LUT_sin[370] = 16'd483;
    LUT_sin[371] = 16'd417;
    LUT_sin[372] = 16'd355;
    LUT_sin[373] = 16'd299;
    LUT_sin[374] = 16'd247;
    LUT_sin[375] = 16'd200;
    LUT_sin[376] = 16'd158;
    LUT_sin[377] = 16'd121;
    LUT_sin[378] = 16'd89;
    LUT_sin[379] = 16'd62;
    LUT_sin[380] = 16'd40;
    LUT_sin[381] = 16'd23;
    LUT_sin[382] = 16'd10;
    LUT_sin[383] = 16'd3;
    LUT_sin[384] = 16'd1;
    LUT_sin[385] = 16'd3;
    LUT_sin[386] = 16'd10;
    LUT_sin[387] = 16'd23;
    LUT_sin[388] = 16'd40;
    LUT_sin[389] = 16'd62;
    LUT_sin[390] = 16'd89;
    LUT_sin[391] = 16'd121;
    LUT_sin[392] = 16'd158;
    LUT_sin[393] = 16'd200;
    LUT_sin[394] = 16'd247;
    LUT_sin[395] = 16'd299;
    LUT_sin[396] = 16'd355;
    LUT_sin[397] = 16'd417;
    LUT_sin[398] = 16'd483;
    LUT_sin[399] = 16'd554;
    LUT_sin[400] = 16'd630;
    LUT_sin[401] = 16'd711;
    LUT_sin[402] = 16'd797;
    LUT_sin[403] = 16'd887;
    LUT_sin[404] = 16'd982;
    LUT_sin[405] = 16'd1083;
    LUT_sin[406] = 16'd1187;
    LUT_sin[407] = 16'd1297;
    LUT_sin[408] = 16'd1411;
    LUT_sin[409] = 16'd1531;
    LUT_sin[410] = 16'd1654;
    LUT_sin[411] = 16'd1783;
    LUT_sin[412] = 16'd1916;
    LUT_sin[413] = 16'd2054;
    LUT_sin[414] = 16'd2196;
    LUT_sin[415] = 16'd2343;
    LUT_sin[416] = 16'd2495;
    LUT_sin[417] = 16'd2651;
    LUT_sin[418] = 16'd2812;
    LUT_sin[419] = 16'd2977;
    LUT_sin[420] = 16'd3146;
    LUT_sin[421] = 16'd3321;
    LUT_sin[422] = 16'd3499;
    LUT_sin[423] = 16'd3682;
    LUT_sin[424] = 16'd3870;
    LUT_sin[425] = 16'd4061;
    LUT_sin[426] = 16'd4257;
    LUT_sin[427] = 16'd4458;
    LUT_sin[428] = 16'd4662;
    LUT_sin[429] = 16'd4871;
    LUT_sin[430] = 16'd5084;
    LUT_sin[431] = 16'd5301;
    LUT_sin[432] = 16'd5523;
    LUT_sin[433] = 16'd5748;
    LUT_sin[434] = 16'd5978;
    LUT_sin[435] = 16'd6211;
    LUT_sin[436] = 16'd6449;
    LUT_sin[437] = 16'd6690;
    LUT_sin[438] = 16'd6936;
    LUT_sin[439] = 16'd7185;
    LUT_sin[440] = 16'd7438;
    LUT_sin[441] = 16'd7695;
    LUT_sin[442] = 16'd7956;
    LUT_sin[443] = 16'd8221;
    LUT_sin[444] = 16'd8489;
    LUT_sin[445] = 16'd8761;
    LUT_sin[446] = 16'd9036;
    LUT_sin[447] = 16'd9315;
    LUT_sin[448] = 16'd9598;
    LUT_sin[449] = 16'd9884;
    LUT_sin[450] = 16'd10173;
    LUT_sin[451] = 16'd10466;
    LUT_sin[452] = 16'd10763;
    LUT_sin[453] = 16'd11062;
    LUT_sin[454] = 16'd11365;
    LUT_sin[455] = 16'd11671;
    LUT_sin[456] = 16'd11980;
    LUT_sin[457] = 16'd12293;
    LUT_sin[458] = 16'd12608;
    LUT_sin[459] = 16'd12927;
    LUT_sin[460] = 16'd13248;
    LUT_sin[461] = 16'd13573;
    LUT_sin[462] = 16'd13900;
    LUT_sin[463] = 16'd14230;
    LUT_sin[464] = 16'd14563;
    LUT_sin[465] = 16'd14899;
    LUT_sin[466] = 16'd15237;
    LUT_sin[467] = 16'd15578;
    LUT_sin[468] = 16'd15922;
    LUT_sin[469] = 16'd16268;
    LUT_sin[470] = 16'd16617;
    LUT_sin[471] = 16'd16968;
    LUT_sin[472] = 16'd17321;
    LUT_sin[473] = 16'd17677;
    LUT_sin[474] = 16'd18035;
    LUT_sin[475] = 16'd18395;
    LUT_sin[476] = 16'd18758;
    LUT_sin[477] = 16'd19122;
    LUT_sin[478] = 16'd19489;
    LUT_sin[479] = 16'd19858;
    LUT_sin[480] = 16'd20228;
    LUT_sin[481] = 16'd20601;
    LUT_sin[482] = 16'd20975;
    LUT_sin[483] = 16'd21351;
    LUT_sin[484] = 16'd21729;
    LUT_sin[485] = 16'd22108;
    LUT_sin[486] = 16'd22489;
    LUT_sin[487] = 16'd22872;
    LUT_sin[488] = 16'd23256;
    LUT_sin[489] = 16'd23641;
    LUT_sin[490] = 16'd24028;
    LUT_sin[491] = 16'd24416;
    LUT_sin[492] = 16'd24806;
    LUT_sin[493] = 16'd25196;
    LUT_sin[494] = 16'd25588;
    LUT_sin[495] = 16'd25981;
    LUT_sin[496] = 16'd26375;
    LUT_sin[497] = 16'd26770;
    LUT_sin[498] = 16'd27166;
    LUT_sin[499] = 16'd27562;
    LUT_sin[500] = 16'd27960;
    LUT_sin[501] = 16'd28358;
    LUT_sin[502] = 16'd28756;
    LUT_sin[503] = 16'd29156;
    LUT_sin[504] = 16'd29556;
    LUT_sin[505] = 16'd29956;
    LUT_sin[506] = 16'd30357;
    LUT_sin[507] = 16'd30758;
    LUT_sin[508] = 16'd31160;
    LUT_sin[509] = 16'd31561;
    LUT_sin[510] = 16'd31963;
    LUT_sin[511] = 16'd32365;
end	
