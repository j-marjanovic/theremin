///////////////////////////////////////////////////////////////////////////////
//   __  __          _____      _         _   _  ______      _______ _____   //
//  |  \/  |   /\   |  __ \    | |  /\   | \ | |/ __ \ \    / /_   _/ ____|  //
//  | \  / |  /  \  | |__) |   | | /  \  |  \| | |  | \ \  / /  | || |       //
//  | |\/| | / /\ \ |  _  /_   | |/ /\ \ | . ` | |  | |\ \/ /   | || |       //
//  | |  | |/ ____ \| | \ \ |__| / ____ \| |\  | |__| | \  /   _| || |____   //
//  |_|  |_/_/    \_\_|  \_\____/_/    \_\_| \_|\____/   \/   |_____\_____|  //
//                                                                           //
//                          JAN MARJANOVIC, 2014                             //
//                                                                           //
///////////////////////////////////////////////////////////////////////////////

`timescale 1ns/100ps

module AD5660_SPI_tb;

localparam Tclk = 20;

//=============================================================================
// Clock
logic clk = 0;
always #(Tclk/2) clk <= !clk;

//=============================================================================
// Reset
logic reset_n=1;
initial begin
	reset_n <= 1;
	#(10*Tclk);
	reset_n <= 0;
	#(10*Tclk);
	reset_n <= 1;
end

//=============================================================================
// Module
localparam BITS = 24;
logic	[BITS-1:0]	in = 24'h85ABCD;
logic				go;
wire				SS_n;
wire				SCLK;	
wire				SDO;

AD5660_SPI #( 
	.BITS	( BITS	) 
) AD5660_SPI_inst ( .* );


//=============================================================================
// Test procedure

initial begin
	$display("========================================");
	$display("=   AD5660_SPI module test procedure   =");
	$display("========================================");

	wait(reset_n == 0);
	$display("%t: Going into reset", $time());

	wait(reset_n == 1);
	$display("%t: Going out of reset", $time());

	#(10*Tclk);
	
	@(posedge clk)
		go	<= 1;

	@(posedge clk)
		go	<= 0;
end

endmodule
